module led_matrix(
    input reg row_data, // inputs a specific row's information
    input 
)